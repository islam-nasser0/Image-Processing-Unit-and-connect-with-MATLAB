module xor_gate (
output c
input a,b,
);
assign c=a^b;
    
endmodule